module ivl_uvm_top;

  `UVM_TESTNAME uvm_test_top;

  initial begin : m_top
    uvm_test_top = new();

  end : m_top
endmodule : ivl_uvm_top

