typedef enum {IDLE, APB_WRITE, APB_READ} kind_e;

