`include "apb_if.sv"
`include "apb_mst_driver.sv"
