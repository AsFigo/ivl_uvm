package apb_pkg;
  import ivl_uvm_pkg::*;
  `include "apb_types.svh"
  `include "apb_mst_xactn.svh"
endpackage : apb_pkg

